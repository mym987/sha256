module sha256_const(addr, k);
  input wire [5:0] addr;
  output wire [31:0] k;

endmodule